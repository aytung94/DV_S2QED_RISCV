
module qed_module(
    input reg [31:0] cpu0_inst,
    input reg [31:0] cpu1_inst
);

endmodule
